interface intf();
  
  logic en;
  logic rst_n;
  logic [2:0] reset_duration;
  logic [2:0] gray_code;
  logic [2:0] count;
  
  
endinterface